module VGA(
    input  wire        PCLK,
    input  wire [7:0]  PRAM,
    output wire        FSYNC,
    output wire        HSYNC,
    output wire        VSYNC,
    output wire        HBLANK,
    output wire        VBLANK,
    output wire [11:0] RGB444
);
    /* horizontal timing parameters */
    localparam H_SYNC  = 95;
    localparam H_BACK  = 143;
    localparam H_DISP  = 783;
    localparam H_FRONT = 799;

    /* vertical timing parameters */
    localparam V_SYNC  = 1;
    localparam V_BACK  = 34;
    localparam V_DISP  = 514;
    localparam V_FRONT = 524;

    /* VGA signal registers */
    reg [9:0]  hcnt = 0;
    reg [9:0]  vcnt = 0;
    reg [11:0] pbuf = 0;

    /* blanking signals */
    assign HBLANK = hcnt > H_DISP || hcnt <= H_BACK;
    assign VBLANK = vcnt > V_DISP || vcnt <= V_BACK;

    /* VGA sync & color signals */
    assign HSYNC        = hcnt > H_SYNC;
    assign VSYNC        = vcnt > V_SYNC;
    assign FSYNC        = vcnt != V_SYNC;
    assign RGB444[11:0] = HBLANK || VBLANK ? 0 : pbuf[11:0];

    /* horizontal timing */
    always @(posedge PCLK) begin
        hcnt <= hcnt == H_FRONT ? 0 : hcnt + 1;
    end

    /* vertical timing */
    always @(posedge PCLK) begin
        if (hcnt == H_FRONT) begin
            vcnt <= vcnt == V_FRONT ? 0 : vcnt + 1;
        end
    end

    /* 256-color mapping */
    always @(PRAM) begin
        case (PRAM)
            8'b00000000: pbuf <= 12'b000000000000;
            8'b00000001: pbuf <= 12'b100000000000;
            8'b00000010: pbuf <= 12'b000010000000;
            8'b00000011: pbuf <= 12'b100010000000;
            8'b00000100: pbuf <= 12'b000000001000;
            8'b00000101: pbuf <= 12'b100000001000;
            8'b00000110: pbuf <= 12'b000010001000;
            8'b00000111: pbuf <= 12'b110011001100;
            8'b00001000: pbuf <= 12'b100010001000;
            8'b00001001: pbuf <= 12'b111100000000;
            8'b00001010: pbuf <= 12'b000011110000;
            8'b00001011: pbuf <= 12'b111111110000;
            8'b00001100: pbuf <= 12'b000000001111;
            8'b00001101: pbuf <= 12'b111100001111;
            8'b00001110: pbuf <= 12'b000011111111;
            8'b00001111: pbuf <= 12'b111111111111;
            8'b00010000: pbuf <= 12'b000000000000;
            8'b00010001: pbuf <= 12'b000000000110;
            8'b00010010: pbuf <= 12'b000000001000;
            8'b00010011: pbuf <= 12'b000000001011;
            8'b00010100: pbuf <= 12'b000000001101;
            8'b00010101: pbuf <= 12'b000000001111;
            8'b00010110: pbuf <= 12'b000001100000;
            8'b00010111: pbuf <= 12'b000001100110;
            8'b00011000: pbuf <= 12'b000001101000;
            8'b00011001: pbuf <= 12'b000001101011;
            8'b00011010: pbuf <= 12'b000001101101;
            8'b00011011: pbuf <= 12'b000001101111;
            8'b00011100: pbuf <= 12'b000010000000;
            8'b00011101: pbuf <= 12'b000010000110;
            8'b00011110: pbuf <= 12'b000010001000;
            8'b00011111: pbuf <= 12'b000010001011;
            8'b00100000: pbuf <= 12'b000010001101;
            8'b00100001: pbuf <= 12'b000010001111;
            8'b00100010: pbuf <= 12'b000010110000;
            8'b00100011: pbuf <= 12'b000010110110;
            8'b00100100: pbuf <= 12'b000010111000;
            8'b00100101: pbuf <= 12'b000010111011;
            8'b00100110: pbuf <= 12'b000010111101;
            8'b00100111: pbuf <= 12'b000010111111;
            8'b00101000: pbuf <= 12'b000011010000;
            8'b00101001: pbuf <= 12'b000011010110;
            8'b00101010: pbuf <= 12'b000011011000;
            8'b00101011: pbuf <= 12'b000011011011;
            8'b00101100: pbuf <= 12'b000011011101;
            8'b00101101: pbuf <= 12'b000011011111;
            8'b00101110: pbuf <= 12'b000011110000;
            8'b00101111: pbuf <= 12'b000011110110;
            8'b00110000: pbuf <= 12'b000011111000;
            8'b00110001: pbuf <= 12'b000011111011;
            8'b00110010: pbuf <= 12'b000011111101;
            8'b00110011: pbuf <= 12'b000011111111;
            8'b00110100: pbuf <= 12'b011000000000;
            8'b00110101: pbuf <= 12'b011000000110;
            8'b00110110: pbuf <= 12'b011000001000;
            8'b00110111: pbuf <= 12'b011000001011;
            8'b00111000: pbuf <= 12'b011000001101;
            8'b00111001: pbuf <= 12'b011000001111;
            8'b00111010: pbuf <= 12'b011001100000;
            8'b00111011: pbuf <= 12'b011001100110;
            8'b00111100: pbuf <= 12'b011001101000;
            8'b00111101: pbuf <= 12'b011001101011;
            8'b00111110: pbuf <= 12'b011001101101;
            8'b00111111: pbuf <= 12'b011001101111;
            8'b01000000: pbuf <= 12'b011010000000;
            8'b01000001: pbuf <= 12'b011010000110;
            8'b01000010: pbuf <= 12'b011010001000;
            8'b01000011: pbuf <= 12'b011010001011;
            8'b01000100: pbuf <= 12'b011010001101;
            8'b01000101: pbuf <= 12'b011010001111;
            8'b01000110: pbuf <= 12'b011010110000;
            8'b01000111: pbuf <= 12'b011010110110;
            8'b01001000: pbuf <= 12'b011010111000;
            8'b01001001: pbuf <= 12'b011010111011;
            8'b01001010: pbuf <= 12'b011010111101;
            8'b01001011: pbuf <= 12'b011010111111;
            8'b01001100: pbuf <= 12'b011011010000;
            8'b01001101: pbuf <= 12'b011011010110;
            8'b01001110: pbuf <= 12'b011011011000;
            8'b01001111: pbuf <= 12'b011011011011;
            8'b01010000: pbuf <= 12'b011011011101;
            8'b01010001: pbuf <= 12'b011011011111;
            8'b01010010: pbuf <= 12'b011011110000;
            8'b01010011: pbuf <= 12'b011011110110;
            8'b01010100: pbuf <= 12'b011011111000;
            8'b01010101: pbuf <= 12'b011011111011;
            8'b01010110: pbuf <= 12'b011011111101;
            8'b01010111: pbuf <= 12'b011011111111;
            8'b01011000: pbuf <= 12'b100000000000;
            8'b01011001: pbuf <= 12'b100000000110;
            8'b01011010: pbuf <= 12'b100000001000;
            8'b01011011: pbuf <= 12'b100000001011;
            8'b01011100: pbuf <= 12'b100000001101;
            8'b01011101: pbuf <= 12'b100000001111;
            8'b01011110: pbuf <= 12'b100001100000;
            8'b01011111: pbuf <= 12'b100001100110;
            8'b01100000: pbuf <= 12'b100001101000;
            8'b01100001: pbuf <= 12'b100001101011;
            8'b01100010: pbuf <= 12'b100001101101;
            8'b01100011: pbuf <= 12'b100001101111;
            8'b01100100: pbuf <= 12'b100010000000;
            8'b01100101: pbuf <= 12'b100010000110;
            8'b01100110: pbuf <= 12'b100010001000;
            8'b01100111: pbuf <= 12'b100010001011;
            8'b01101000: pbuf <= 12'b100010001101;
            8'b01101001: pbuf <= 12'b100010001111;
            8'b01101010: pbuf <= 12'b100010110000;
            8'b01101011: pbuf <= 12'b100010110110;
            8'b01101100: pbuf <= 12'b100010111000;
            8'b01101101: pbuf <= 12'b100010111011;
            8'b01101110: pbuf <= 12'b100010111101;
            8'b01101111: pbuf <= 12'b100010111111;
            8'b01110000: pbuf <= 12'b100011010000;
            8'b01110001: pbuf <= 12'b100011010110;
            8'b01110010: pbuf <= 12'b100011011000;
            8'b01110011: pbuf <= 12'b100011011011;
            8'b01110100: pbuf <= 12'b100011011101;
            8'b01110101: pbuf <= 12'b100011011111;
            8'b01110110: pbuf <= 12'b100011110000;
            8'b01110111: pbuf <= 12'b100011110110;
            8'b01111000: pbuf <= 12'b100011111000;
            8'b01111001: pbuf <= 12'b100011111011;
            8'b01111010: pbuf <= 12'b100011111101;
            8'b01111011: pbuf <= 12'b100011111111;
            8'b01111100: pbuf <= 12'b101100000000;
            8'b01111101: pbuf <= 12'b101100000110;
            8'b01111110: pbuf <= 12'b101100001000;
            8'b01111111: pbuf <= 12'b101100001011;
            8'b10000000: pbuf <= 12'b101100001101;
            8'b10000001: pbuf <= 12'b101100001111;
            8'b10000010: pbuf <= 12'b101101100000;
            8'b10000011: pbuf <= 12'b101101100110;
            8'b10000100: pbuf <= 12'b101101101000;
            8'b10000101: pbuf <= 12'b101101101011;
            8'b10000110: pbuf <= 12'b101101101101;
            8'b10000111: pbuf <= 12'b101101101111;
            8'b10001000: pbuf <= 12'b101110000000;
            8'b10001001: pbuf <= 12'b101110000110;
            8'b10001010: pbuf <= 12'b101110001000;
            8'b10001011: pbuf <= 12'b101110001011;
            8'b10001100: pbuf <= 12'b101110001101;
            8'b10001101: pbuf <= 12'b101110001111;
            8'b10001110: pbuf <= 12'b101110110000;
            8'b10001111: pbuf <= 12'b101110110110;
            8'b10010000: pbuf <= 12'b101110111000;
            8'b10010001: pbuf <= 12'b101110111011;
            8'b10010010: pbuf <= 12'b101110111101;
            8'b10010011: pbuf <= 12'b101110111111;
            8'b10010100: pbuf <= 12'b101111010000;
            8'b10010101: pbuf <= 12'b101111010110;
            8'b10010110: pbuf <= 12'b101111011000;
            8'b10010111: pbuf <= 12'b101111011011;
            8'b10011000: pbuf <= 12'b101111011101;
            8'b10011001: pbuf <= 12'b101111011111;
            8'b10011010: pbuf <= 12'b101111110000;
            8'b10011011: pbuf <= 12'b101111110110;
            8'b10011100: pbuf <= 12'b101111111000;
            8'b10011101: pbuf <= 12'b101111111011;
            8'b10011110: pbuf <= 12'b101111111101;
            8'b10011111: pbuf <= 12'b101111111111;
            8'b10100000: pbuf <= 12'b110100000000;
            8'b10100001: pbuf <= 12'b110100000110;
            8'b10100010: pbuf <= 12'b110100001000;
            8'b10100011: pbuf <= 12'b110100001011;
            8'b10100100: pbuf <= 12'b110100001101;
            8'b10100101: pbuf <= 12'b110100001111;
            8'b10100110: pbuf <= 12'b110101100000;
            8'b10100111: pbuf <= 12'b110101100110;
            8'b10101000: pbuf <= 12'b110101101000;
            8'b10101001: pbuf <= 12'b110101101011;
            8'b10101010: pbuf <= 12'b110101101101;
            8'b10101011: pbuf <= 12'b110101101111;
            8'b10101100: pbuf <= 12'b110110000000;
            8'b10101101: pbuf <= 12'b110110000110;
            8'b10101110: pbuf <= 12'b110110001000;
            8'b10101111: pbuf <= 12'b110110001011;
            8'b10110000: pbuf <= 12'b110110001101;
            8'b10110001: pbuf <= 12'b110110001111;
            8'b10110010: pbuf <= 12'b110110110000;
            8'b10110011: pbuf <= 12'b110110110110;
            8'b10110100: pbuf <= 12'b110110111000;
            8'b10110101: pbuf <= 12'b110110111011;
            8'b10110110: pbuf <= 12'b110110111101;
            8'b10110111: pbuf <= 12'b110110111111;
            8'b10111000: pbuf <= 12'b110111010000;
            8'b10111001: pbuf <= 12'b110111010110;
            8'b10111010: pbuf <= 12'b110111011000;
            8'b10111011: pbuf <= 12'b110111011011;
            8'b10111100: pbuf <= 12'b110111011101;
            8'b10111101: pbuf <= 12'b110111011111;
            8'b10111110: pbuf <= 12'b110111110000;
            8'b10111111: pbuf <= 12'b110111110110;
            8'b11000000: pbuf <= 12'b110111111000;
            8'b11000001: pbuf <= 12'b110111111011;
            8'b11000010: pbuf <= 12'b110111111101;
            8'b11000011: pbuf <= 12'b110111111111;
            8'b11000100: pbuf <= 12'b111100000000;
            8'b11000101: pbuf <= 12'b111100000110;
            8'b11000110: pbuf <= 12'b111100001000;
            8'b11000111: pbuf <= 12'b111100001011;
            8'b11001000: pbuf <= 12'b111100001101;
            8'b11001001: pbuf <= 12'b111100001111;
            8'b11001010: pbuf <= 12'b111101100000;
            8'b11001011: pbuf <= 12'b111101100110;
            8'b11001100: pbuf <= 12'b111101101000;
            8'b11001101: pbuf <= 12'b111101101011;
            8'b11001110: pbuf <= 12'b111101101101;
            8'b11001111: pbuf <= 12'b111101101111;
            8'b11010000: pbuf <= 12'b111110000000;
            8'b11010001: pbuf <= 12'b111110000110;
            8'b11010010: pbuf <= 12'b111110001000;
            8'b11010011: pbuf <= 12'b111110001011;
            8'b11010100: pbuf <= 12'b111110001101;
            8'b11010101: pbuf <= 12'b111110001111;
            8'b11010110: pbuf <= 12'b111110110000;
            8'b11010111: pbuf <= 12'b111110110110;
            8'b11011000: pbuf <= 12'b111110111000;
            8'b11011001: pbuf <= 12'b111110111011;
            8'b11011010: pbuf <= 12'b111110111101;
            8'b11011011: pbuf <= 12'b111110111111;
            8'b11011100: pbuf <= 12'b111111010000;
            8'b11011101: pbuf <= 12'b111111010110;
            8'b11011110: pbuf <= 12'b111111011000;
            8'b11011111: pbuf <= 12'b111111011011;
            8'b11100000: pbuf <= 12'b111111011101;
            8'b11100001: pbuf <= 12'b111111011111;
            8'b11100010: pbuf <= 12'b111111110000;
            8'b11100011: pbuf <= 12'b111111110110;
            8'b11100100: pbuf <= 12'b111111111000;
            8'b11100101: pbuf <= 12'b111111111011;
            8'b11100110: pbuf <= 12'b111111111101;
            8'b11100111: pbuf <= 12'b111111111111;
            8'b11101000: pbuf <= 12'b000100010001;
            8'b11101001: pbuf <= 12'b001000100010;
            8'b11101010: pbuf <= 12'b001000100010;
            8'b11101011: pbuf <= 12'b001100110011;
            8'b11101100: pbuf <= 12'b001100110011;
            8'b11101101: pbuf <= 12'b010001000100;
            8'b11101110: pbuf <= 12'b010001000100;
            8'b11101111: pbuf <= 12'b010101010101;
            8'b11110000: pbuf <= 12'b011001100110;
            8'b11110001: pbuf <= 12'b011001100110;
            8'b11110010: pbuf <= 12'b011101110111;
            8'b11110011: pbuf <= 12'b011101110111;
            8'b11110100: pbuf <= 12'b100010001000;
            8'b11110101: pbuf <= 12'b100110011001;
            8'b11110110: pbuf <= 12'b100110011001;
            8'b11110111: pbuf <= 12'b101010101010;
            8'b11111000: pbuf <= 12'b101010101010;
            8'b11111001: pbuf <= 12'b101110111011;
            8'b11111010: pbuf <= 12'b110011001100;
            8'b11111011: pbuf <= 12'b110011001100;
            8'b11111100: pbuf <= 12'b110111011101;
            8'b11111101: pbuf <= 12'b110111011101;
            8'b11111110: pbuf <= 12'b111011101110;
            8'b11111111: pbuf <= 12'b111011101110;
        endcase
    end
endmodule

module main(
    input  wire clk,
    // input  wire P1_1,
    // input  wire P1_2,
    // input  wire P1_3,
    // input  wire P1_4,
    // input  wire P1_9,
    // input  wire P1_10,
    // input  wire P1_11,
    // input  wire P1_12,
    output wire P2_1,
    output wire P2_2,
    output wire P2_3,
    output wire P2_4,
    output wire P2_9,
    output wire P2_10,
    output wire P2_11,
    output wire P2_12,
    output wire P3_1,
    output wire P3_2,
    output wire P3_9,
    output wire P3_10,
    output wire P3_11,
    output wire P3_12,
    output wire P4_1,
    output wire P4_2
);
    wire pclk;
    wire locked;

    /* pixel clock @ 25.125MHz */
    PLL pll(
        .clock_in  (clk),
        .clock_out (pclk),
        .locked    (locked)
    );

    /* sync & blanking signals */
    wire fsync;
    wire hsync;
    wire vsync;
    wire hblank;
    wire vblank;

    /* connect the sync signals */
    assign P3_1 = hsync;
    assign P3_2 = vsync;

    /* frame sync & pixel clock */
    assign P4_1 = fsync;
    assign P4_2 = hblank | vblank | ~pclk;

    /* connect the color signals */
    // wire [7:0] pixel = {
    //     P1_12,
    //     P1_11,
    //     P1_10,
    //     P1_9,
    //     P1_1,
    //     P1_2,
    //     P1_3,
    //     P1_4
    // };

    reg [5:0] col = 0;
    reg [9:0] cnt = 0;
    reg [7:0] pixel = 0;
    always @(posedge pclk) begin
        if (~fsync) begin
            col <= 0;
            cnt <= 0;
            pixel <= 0;
        end else if (~hblank && ~vblank) begin
            if (col != 39) begin
                col <= col + 1;
            end else begin
                col <= 0;
                if (cnt == 479) begin
                    cnt   <= 0;
                    pixel <= pixel + 1;
                end else if (cnt[3:0] != 4'b1111) begin
                    cnt   <= cnt + 1;
                    pixel <= pixel + 1;
                end else begin
                    cnt   <= cnt + 1;
                    pixel <= pixel - 15;
                end
            end
        end
    end

    /* VGA module */
    VGA vga(
        .PCLK   (pclk),
        .PRAM   (pixel),
        .FSYNC  (fsync),
        .HSYNC  (hsync),
        .VSYNC  (vsync),
        .HBLANK (hblank),
        .VBLANK (vblank),
        .RGB444 ({P2_9, P2_10, P2_11, P2_12, P3_9, P3_10, P3_11, P3_12, P2_4, P2_3, P2_2, P2_1})
    );
endmodule
